Library IEEE;
use IEEE.std_logic_1164.all;

--Entity
Entity  is
port(
A:in STD_LOGIC;
B:in STD_LOGIC;
Cin:in STD_LOGIC;
C0,sum:out STD_LOGIC
);

architecture